

module dummy_dut;
endmodule
