//------------------------------------------------------------------------------
//File       : dummy_dut.sv
//Author     : Krishna Gupta/1BM23EC123
//Created    : 2026-01-29
//Module     : dummy_dut
//Project    : SystemVerilog and Verification (23EC6PE2SV)
//Faculty    : Prof. Ajaykumar Devarapalli
//Description: A placeholder dummy DUT for the class-based Packet verification lab.
//------------------------------------------------------------------------------

module dummy_dut;
endmodule
